package MemoryPkg;

  import ROM::*;
  export ROM::*;

endpackage