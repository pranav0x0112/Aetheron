package TileLinkPkg;

  import TLMasterXactor::*;
  import TLSlaveXactor::*;
  import TLTypes::*;

  export TLMasterXactorIfc;
  export TLSlaveXactorIfc;
  export TLTypes::*;

endpackage