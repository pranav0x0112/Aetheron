package PeripheralsPkg;

  import GPIO::*;

  export GPIO::*;

endpackage