package TileLinkPkg;

  import TLMasterXactor::*;
  import TLSlaveXactor::*;
  import TLTypes::*;

  export TLMasterXactor::*;
  export TLSlaveXactor::*;
  export TLTypes::*;

endpackage